module ALUcontroller (ports);
    
endmodule
